`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/02/2020 02:04:14 PM
// Design Name: 
// Module Name: tb_multiplier
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_multiplier( );
    parameter N=16,M=4;
    reg [N-1:0] A,B;
    wire [2*N-1:0] PRODUCT;
    
    MAIN_1 #(N,M) m1  (A,B,PRODUCT);
    
    //Testing using random inputs
    initial begin
//    A = 8'b11111111; B = 8'b10001000; #10
//    A = 8'b11111111; B = 8'b10001001; #10
//    A = 8'b11111111; B = 8'b11111111; #10
//    B = 8'b10011011; A = 8'b10100111; #10
    
    A = 16'b1111111111111111; B = 16'b1000100010001000; #10
    A = 16'b1111111111111111; B = 16'b1000100111111111; #10
    A = 16'b1111111111111111; B = 16'b1111111111111111; #10
    B = 16'b1001101110011011; A = 16'b1010011110100111; #10
    
//    A = 32'b11111111111111111111111111111111; B = 32'b10001000100010001000100010001000; #10
//    A = 32'b11111111111111111000100010001000; B = 32'b10001001111111111000100010001000; #10
//    A = 32'b11111111111111111000100010001000; B = 32'b11111111111111111000100010001000; #10
//    B = 32'b10011011100110111000100010001000; A = 32'b10100111101001111000100010001000; #10
    
    $finish;
    end
endmodule
